module kooft(input a, output b);

endmodule
